library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity EntidadControlAscensor is
    Port ( PisoVoy : in  STD_LOGIC_VECTOR (3 downto 0);
           PisoEstoy : in  STD_LOGIC_VECTOR (3 downto 0);
           ControlMotor : out  STD_LOGIC_VECTOR (1 downto 0)
			  );
end EntidadControlAscensor;

architecture Behavioral of EntidadControlAscensor is


	component DecodificadorBinarioEntero 
	port (
			EntradaBinaria: in std_logic_vector (3 downto 0);
			SalidaEntera : out  INTEGER
			);
	end component;

	component Comparador
	port (
			PisoVoy: in INTEGER;
			PisoEstoy: in INTEGER;
			ControlMotor : out  STD_LOGIC_VECTOR (1 downto 0)
			);
	end component;
	
	--signal declaration
	signal SigPisoVoy, SigPisoEstoy : INTEGER;
	
begin

	Inst_decodificadorVoy: DecodificadorBinarioEntero port map (
		EntradaBinaria => PisoVoy, 
		SalidaEntera => SigPisoVoy  	
	);

	Inst_decodificadorEstoy: DecodificadorBinarioEntero port map (
		EntradaBinaria => PisoEstoy, 
		SalidaEntera => SigPisoEstoy
	);
	
	Inst_Comparador: Comparador port map (
		PisoVoy => SigPisoVoy,
		PisoEstoy => SigPisoEstoy, 	
		ControlMotor => ControlMotor
	);

end Behavioral;